`timescale 1ns / 1ps


module Ctr(
    input [5:0] opCode,


    output reg regDest,
    output reg aluSrc,
    output reg memToReg,
    output reg regWrite,
    output reg memRead,
    output reg memWrite,
    output reg Branch,
    output reg [2:0] ALUop,
    output reg Jump,
    output reg jumpTarget,
    output reg Call,
    output reg [1:0] Signed,
    output reg branchEqual
    );
    always @(opCode)
    begin
        case(opCode)
            6'b000000://add,addu,sub,subu,and,or,xor,nor,slt,jr,sltu,sll,srl,sra,sllv,srlv,srav,jr
            begin
                regDest=1;
                aluSrc=0;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b010;
                Signed=0;
            end
            6'b000010://jump
            begin
                regDest=0;
                aluSrc=0;
                memToReg=0;
                regWrite=0;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=1;
                jumpTarget=1;
                Call=0;
                ALUop=3'b000;
                Signed=0;
            end
            6'b000011://jal
            begin
                regDest=1;
                aluSrc=0;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=1;
                jumpTarget=1;
                Call=1;
                ALUop=3'b000;
                Signed=0;
            end
            6'b001000://addi
            begin
                regDest=0;
                aluSrc=1;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b000;
                Signed=0;
            end
            6'b001001://addiu
            begin
                regDest=0;
                aluSrc=1;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b000;
                Signed=1;
            end 
            6'b001100://andi
            begin
                regDest=0;
                aluSrc=1;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b000;
                Signed=0;
            end
            6'b001101://ori
            begin
                regDest=0;
                aluSrc=1;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b000;
                Signed=0;
            end
            6'b001110://xori
            begin
                regDest=0;
                aluSrc=1;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b000;
                Signed=0;
            end
            6'b001111://lui
            begin
                regDest=0;
                aluSrc=1;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b000;
                Signed=2'b10;
            end
            6'b100011://lw
            begin
                regDest=0;
                aluSrc=1;
                memToReg=1;
                regWrite=1;
                memRead=1;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b000;
                Signed=1;
            end
            6'b101011://sw
            begin
                regDest=1;
                aluSrc=1;
                memToReg=0;
                regWrite=0;
                memRead=0;
                memWrite=1;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b000;
                Signed=1;
            end
            6'b000100://beq
            begin
                regDest=1;
                aluSrc=0;
                regWrite=0;
                memToReg=0;
                memRead=0;
                memWrite=0;
                Branch=1;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b001;
                Signed=1;
                branchEqual=1;
            end
            6'b000101://bne
            begin
                regDest=1;
                aluSrc=0;
                regWrite=0;
                memToReg=0;
                memRead=0;
                memWrite=0;
                Branch=1;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b001;
                Signed=1;
                branchEqual=0;
            end
            6'b001010://slti
            begin
                regDest=0;
                aluSrc=1;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b111;
                Signed=1;
            end
            6'b001011://sltiu
            begin
                regDest=0;
                aluSrc=1;
                memToReg=0;
                regWrite=1;
                memRead=0;
                memWrite=0;
                Branch=0;
                Jump=0;
                jumpTarget=0;
                Call=0;
                ALUop=3'b010;
                Signed=0;
            end    
        endcase
    end
endmodule
